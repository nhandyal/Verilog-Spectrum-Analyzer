`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    23:01:29 04/30/2012 
// Design Name: 
// Module Name:    complexMult_TopBranch 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module complexMultN(DinAR, DinAI, DinBR, DinBI, DoutR, DoutI);

	input 	[17:0] DinAR, DinAI, DinBR, DinBI;
	output 	[17:0] DoutR, DoutI;
	
	


endmodule
